** Profile: "SCHEMATIC1-example2"  [ C:\Users\Huang Xianmin\Desktop\Pspice_simulation_file\test-PSpiceFiles\SCHEMATIC1\example2.sim ] 

** Creating circuit file "example2.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of D:\Cadence\SPB_16.5\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V1 0v 5v 1v 
.TEMP 20 100 200
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
