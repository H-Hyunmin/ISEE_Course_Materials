module decrement (
    input [7:0] A,
    output [7:0] F
);
    assign F = A - 1;
endmodule