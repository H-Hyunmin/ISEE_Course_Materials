module increment (
    input [3:0] A,
    output [3:0] F
);
    assign F = A + 1;
    
endmodule